`include "cpu_ram_if.vh"
`timescale 1 ns / 1 ns

