`ifndef ICACHE_PKG_VH
`define ICACHE_PKG_VH
package icache_pkg;

  typedef logic [26:0] tags;

endpackage
`endif //ICACHE_PKG_VH
